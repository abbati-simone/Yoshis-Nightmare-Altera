parameter ROM_0_messages_len=146;
parameter ROM_0_note_min=67;
parameter ROM_0_note_max=84;
parameter ROM_0_delay_min=0;
parameter ROM_0_delay_max=960;
parameter ROM_0_messages_address_bits=8;
parameter ROM_0_note_nbit=5;
parameter ROM_0_delay_nbit=10;

