parameter ROMS_number=2;
parameter note_max_bits=5;
parameter address_max_bits=12;
parameter delay_max_bits=14;
parameter ticks_per_beat=1024;
parameter BPM=400;
parameter BPS=6.666666666666667;
parameter ticks_hz=6827;
parameter delay_clocks_per_tick=1000;
parameter delay_clock_hz=6827000;
parameter delay_reg_bits=36;

