parameter ROM_0_messages_len=2448;
parameter ROM_0_note_min=55;
parameter ROM_0_note_max=84;
parameter ROM_0_delay_min=0;
parameter ROM_0_delay_max=9213;
parameter ROM_0_messages_address_bits=12;
parameter ROM_0_note_nbit=5;
parameter ROM_0_delay_nbit=14;

