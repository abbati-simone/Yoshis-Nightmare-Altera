parameter ROMS_number=1;
parameter note_max_bits=5;
parameter address_max_bits=8;
parameter delay_max_bits=10;
parameter ticks_per_beat=240;
parameter BPM=120;
parameter BPS=2.0;
parameter ticks_hz=480;
parameter delay_clocks_per_tick=1000;
parameter delay_clock_hz=480000;
parameter delay_reg_bits=29;

