parameter ROM_1_messages_len=1104;
parameter ROM_1_note_min=43;
parameter ROM_1_note_max=65;
parameter ROM_1_delay_min=0;
parameter ROM_1_delay_max=6168;
parameter ROM_1_messages_address_bits=11;
parameter ROM_1_note_nbit=5;
parameter ROM_1_delay_nbit=13;

