module notes_sequence_Yoshi2_0(
	input clk,
	input [8:0] address,
	output reg [4:0] note,
	output reg note_on,
	output reg [11:0] delay
);

reg [17:0] note_;

always @(posedge clk) begin
case(address)
0:note_<=18'b101000000000000000;
1:note_<=18'b001000000011110000;
2:note_<=18'b100111000000000000;
3:note_<=18'b000111000011110000;
4:note_<=18'b101000000000000000;
5:note_<=18'b001000000111100000;
6:note_<=18'b100101000000000000;
7:note_<=18'b000101000111100000;
8:note_<=18'b100101000000000000;
9:note_<=18'b000101001011010000;
10:note_<=18'b100011000000000000;
11:note_<=18'b000011000011110000;
12:note_<=18'b100001000000000000;
13:note_<=18'b000001000111100000;
14:note_<=18'b100101000000000000;
15:note_<=18'b000101000111100000;
16:note_<=18'b100101000000000000;
17:note_<=18'b000101001111000000;
18:note_<=18'b100110000000000000;
19:note_<=18'b000110000011110000;
20:note_<=18'b100110000000000000;
21:note_<=18'b000110000011110000;
22:note_<=18'b100101000011110000;
23:note_<=18'b000101000011110000;
24:note_<=18'b100110000000000000;
25:note_<=18'b000110000111100000;
26:note_<=18'b101000000000000000;
27:note_<=18'b001000000111100000;
28:note_<=18'b101010000000000000;
29:note_<=18'b001010010110100000;
30:note_<=18'b100110000000000000;
31:note_<=18'b000110000011110000;
32:note_<=18'b100101000000000000;
33:note_<=18'b000101000011110000;
34:note_<=18'b100110000000000000;
35:note_<=18'b000110000111100000;
36:note_<=18'b100011000000000000;
37:note_<=18'b000011000111100000;
38:note_<=18'b100011000000000000;
39:note_<=18'b000011001011010000;
40:note_<=18'b100001000000000000;
41:note_<=18'b000001000011110000;
42:note_<=18'b100000000000000000;
43:note_<=18'b000000000111100000;
44:note_<=18'b100011000000000000;
45:note_<=18'b000011000111100000;
46:note_<=18'b100011000000000000;
47:note_<=18'b000011001111000000;
48:note_<=18'b100101000000000000;
49:note_<=18'b000101000011110000;
50:note_<=18'b100101000000000000;
51:note_<=18'b000101000011110000;
52:note_<=18'b100011000011110000;
53:note_<=18'b000011000011110000;
54:note_<=18'b100101000000000000;
55:note_<=18'b000101000111100000;
56:note_<=18'b100011000000000000;
57:note_<=18'b000011000111100000;
58:note_<=18'b100001000000000000;
59:note_<=18'b000001010110100000;
60:note_<=18'b101000000000000000;
61:note_<=18'b001000000011110000;
62:note_<=18'b100111000000000000;
63:note_<=18'b000111000011110000;
64:note_<=18'b101000000000000000;
65:note_<=18'b001000000111100000;
66:note_<=18'b100101000000000000;
67:note_<=18'b000101000111100000;
68:note_<=18'b100101000000000000;
69:note_<=18'b000101001011010000;
70:note_<=18'b100011000000000000;
71:note_<=18'b000011000011110000;
72:note_<=18'b100001000000000000;
73:note_<=18'b000001000111100000;
74:note_<=18'b100101000000000000;
75:note_<=18'b000101000111100000;
76:note_<=18'b100101000000000000;
77:note_<=18'b000101001111000000;
78:note_<=18'b100110000000000000;
79:note_<=18'b000110000011110000;
80:note_<=18'b100110000000000000;
81:note_<=18'b000110000011110000;
82:note_<=18'b100101000011110000;
83:note_<=18'b000101000011110000;
84:note_<=18'b100110000000000000;
85:note_<=18'b000110000111100000;
86:note_<=18'b101000000000000000;
87:note_<=18'b001000000111100000;
88:note_<=18'b101010000000000000;
89:note_<=18'b001010010110100000;
90:note_<=18'b100110000000000000;
91:note_<=18'b000110000011110000;
92:note_<=18'b100101000000000000;
93:note_<=18'b000101000011110000;
94:note_<=18'b100110000000000000;
95:note_<=18'b000110000111100000;
96:note_<=18'b100011000000000000;
97:note_<=18'b000011000111100000;
98:note_<=18'b100011000000000000;
99:note_<=18'b000011001011010000;
100:note_<=18'b100001000000000000;
101:note_<=18'b000001000011110000;
102:note_<=18'b100000000000000000;
103:note_<=18'b000000000111100000;
104:note_<=18'b100011000000000000;
105:note_<=18'b000011000111100000;
106:note_<=18'b100011000000000000;
107:note_<=18'b000011001111000000;
108:note_<=18'b100101000000000000;
109:note_<=18'b000101000011110000;
110:note_<=18'b100101000000000000;
111:note_<=18'b000101000011110000;
112:note_<=18'b100011000011110000;
113:note_<=18'b000011000011110000;
114:note_<=18'b100101000000000000;
115:note_<=18'b000101000111100000;
116:note_<=18'b100011000000000000;
117:note_<=18'b000011000111100000;
118:note_<=18'b100001000000000000;
119:note_<=18'b000001000111100000;
120:note_<=18'b100001000000000000;
121:note_<=18'b000001000111100000;
122:note_<=18'b100011000000000000;
123:note_<=18'b000011000111100000;
124:note_<=18'b100101000000000000;
125:note_<=18'b000101000111100000;
126:note_<=18'b100110000000000000;
127:note_<=18'b000110001111000000;
128:note_<=18'b101010000000000000;
129:note_<=18'b001010010110100000;
130:note_<=18'b101010000000000000;
131:note_<=18'b001010000111100000;
132:note_<=18'b101000000000000000;
133:note_<=18'b001000000111100000;
134:note_<=18'b100110000000000000;
135:note_<=18'b000110000111100000;
136:note_<=18'b100101000000000000;
137:note_<=18'b000101001111000000;
138:note_<=18'b101000000000000000;
139:note_<=18'b001000010110100000;
140:note_<=18'b101000000000000000;
141:note_<=18'b001000000111100000;
142:note_<=18'b100110000000000000;
143:note_<=18'b000110000111100000;
144:note_<=18'b100101000000000000;
145:note_<=18'b000101000111100000;
146:note_<=18'b100011000000000000;
147:note_<=18'b000011001111000000;
148:note_<=18'b100110000000000000;
149:note_<=18'b000110010110100000;
150:note_<=18'b100110000000000000;
151:note_<=18'b000110000111100000;
152:note_<=18'b100101000000000000;
153:note_<=18'b000101000111100000;
154:note_<=18'b100011000000000000;
155:note_<=18'b000011000111100000;
156:note_<=18'b100101000000000000;
157:note_<=18'b000101001111000000;
158:note_<=18'b100110000000000000;
159:note_<=18'b000110001111000000;
160:note_<=18'b101000000000000000;
161:note_<=18'b001000000111100000;
162:note_<=18'b100001000000000000;
163:note_<=18'b000001000111100000;
164:note_<=18'b100011000000000000;
165:note_<=18'b000011000111100000;
166:note_<=18'b100101000000000000;
167:note_<=18'b000101000111100000;
168:note_<=18'b100110000000000000;
169:note_<=18'b000110001111000000;
170:note_<=18'b101010000000000000;
171:note_<=18'b001010010110100000;
172:note_<=18'b101010000000000000;
173:note_<=18'b001010000111100000;
174:note_<=18'b101100000000000000;
175:note_<=18'b001100000111100000;
176:note_<=18'b101101000000000000;
177:note_<=18'b001101000111100000;
178:note_<=18'b110001000000000000;
179:note_<=18'b010001001111000000;
180:note_<=18'b101111000000000000;
181:note_<=18'b001111001111000000;
182:note_<=18'b101110000000000000;
183:note_<=18'b001110001111000000;
184:note_<=18'b101001000000000000;
185:note_<=18'b001001000111100000;
186:note_<=18'b101010000000000000;
187:note_<=18'b001010000111100000;
188:note_<=18'b101111000000000000;
189:note_<=18'b001111001111000000;
190:note_<=18'b101010000000000000;
191:note_<=18'b001010001111000000;
192:note_<=18'b101000000000000000;
193:note_<=18'b001000000111100000;
194:note_<=18'b110001000000000000;
195:note_<=18'b010001000111100000;
196:note_<=18'b101111000000000000;
197:note_<=18'b001111000111100000;
198:note_<=18'b101100000000000000;
199:note_<=18'b001100000111100000;
200:note_<=18'b101101000000000000;
201:note_<=18'b001101110100100000;
202:note_<=18'b101000000000000000;
203:note_<=18'b001000000011110000;
204:note_<=18'b100111000000000000;
205:note_<=18'b000111000011110000;
206:note_<=18'b101000000000000000;
207:note_<=18'b001000000111100000;
208:note_<=18'b100101000000000000;
209:note_<=18'b000101000111100000;
210:note_<=18'b100101000000000000;
211:note_<=18'b000101001011010000;
212:note_<=18'b100011000000000000;
213:note_<=18'b000011000011110000;
214:note_<=18'b100001000000000000;
215:note_<=18'b000001000111100000;
216:note_<=18'b100101000000000000;
217:note_<=18'b000101000111100000;
218:note_<=18'b100101000000000000;
219:note_<=18'b000101001111000000;
220:note_<=18'b100110000000000000;
221:note_<=18'b000110000011110000;
222:note_<=18'b100110000000000000;
223:note_<=18'b000110000011110000;
224:note_<=18'b100101000011110000;
225:note_<=18'b000101000011110000;
226:note_<=18'b100110000000000000;
227:note_<=18'b000110000111100000;
228:note_<=18'b101000000000000000;
229:note_<=18'b001000000111100000;
230:note_<=18'b101010000000000000;
231:note_<=18'b001010010110100000;
232:note_<=18'b100110000000000000;
233:note_<=18'b000110000011110000;
234:note_<=18'b100101000000000000;
235:note_<=18'b000101000011110000;
236:note_<=18'b100110000000000000;
237:note_<=18'b000110000111100000;
238:note_<=18'b100011000000000000;
239:note_<=18'b000011000111100000;
240:note_<=18'b100011000000000000;
241:note_<=18'b000011001011010000;
242:note_<=18'b100001000000000000;
243:note_<=18'b000001000011110000;
244:note_<=18'b100000000000000000;
245:note_<=18'b000000000111100000;
246:note_<=18'b100011000000000000;
247:note_<=18'b000011000111100000;
248:note_<=18'b100011000000000000;
249:note_<=18'b000011001111000000;
250:note_<=18'b100101000000000000;
251:note_<=18'b000101000011110000;
252:note_<=18'b100101000000000000;
253:note_<=18'b000101000011110000;
254:note_<=18'b100011000011110000;
255:note_<=18'b000011000011110000;
256:note_<=18'b100101000000000000;
257:note_<=18'b000101000111100000;
258:note_<=18'b100011000000000000;
259:note_<=18'b000011000111100000;
260:note_<=18'b100001000000000000;
261:note_<=18'b000001010110100000;
262:note_<=18'b101000000000000000;
263:note_<=18'b001000000011110000;
264:note_<=18'b100111000000000000;
265:note_<=18'b000111000011110000;
266:note_<=18'b101000000000000000;
267:note_<=18'b001000000111100000;
268:note_<=18'b100101000000000000;
269:note_<=18'b000101000111100000;
270:note_<=18'b100101000000000000;
271:note_<=18'b000101001011010000;
272:note_<=18'b100011000000000000;
273:note_<=18'b000011000011110000;
274:note_<=18'b100001000000000000;
275:note_<=18'b000001000111100000;
276:note_<=18'b100101000000000000;
277:note_<=18'b000101000111100000;
278:note_<=18'b100101000000000000;
279:note_<=18'b000101001111000000;
280:note_<=18'b100110000000000000;
281:note_<=18'b000110000011110000;
282:note_<=18'b100110000000000000;
283:note_<=18'b000110000011110000;
284:note_<=18'b100101000011110000;
285:note_<=18'b000101000011110000;
286:note_<=18'b100110000000000000;
287:note_<=18'b000110000111100000;
288:note_<=18'b101000000000000000;
289:note_<=18'b001000000111100000;
290:note_<=18'b101010000000000000;
291:note_<=18'b001010010110100000;
292:note_<=18'b100110000000000000;
293:note_<=18'b000110000011110000;
294:note_<=18'b100101000000000000;
295:note_<=18'b000101000011110000;
296:note_<=18'b100110000000000000;
297:note_<=18'b000110000111100000;
298:note_<=18'b100011000000000000;
299:note_<=18'b000011000111100000;
300:note_<=18'b100011000000000000;
301:note_<=18'b000011001011010000;
302:note_<=18'b100001000000000000;
303:note_<=18'b000001000011110000;
304:note_<=18'b100000000000000000;
305:note_<=18'b000000000111100000;
306:note_<=18'b100011000000000000;
307:note_<=18'b000011000111100000;
308:note_<=18'b100011000000000000;
309:note_<=18'b000011001111000000;
310:note_<=18'b100101000000000000;
311:note_<=18'b000101000011110000;
312:note_<=18'b100101000000000000;
313:note_<=18'b000101000011110000;
314:note_<=18'b100011000011110000;
315:note_<=18'b000011000011110000;
316:note_<=18'b100101000000000000;
317:note_<=18'b000101000111100000;
318:note_<=18'b100011000000000000;
319:note_<=18'b000011000111100000;
320:note_<=18'b100001000000000000;
321:note_<=18'b000001000111100000;
322:note_<=18'b100001000000000000;
323:note_<=18'b000001000111100000;
324:note_<=18'b100011000000000000;
325:note_<=18'b000011000111100000;
326:note_<=18'b100101000000000000;
327:note_<=18'b000101000111100000;
328:note_<=18'b100110000000000000;
329:note_<=18'b000110001111000000;
330:note_<=18'b101010000000000000;
331:note_<=18'b001010010110100000;
332:note_<=18'b101010000000000000;
333:note_<=18'b001010000111100000;
334:note_<=18'b101000000000000000;
335:note_<=18'b001000000111100000;
336:note_<=18'b100110000000000000;
337:note_<=18'b000110000111100000;
338:note_<=18'b100101000000000000;
339:note_<=18'b000101001111000000;
340:note_<=18'b101000000000000000;
341:note_<=18'b001000010110100000;
342:note_<=18'b101000000000000000;
343:note_<=18'b001000000111100000;
344:note_<=18'b100110000000000000;
345:note_<=18'b000110000111100000;
346:note_<=18'b100101000000000000;
347:note_<=18'b000101000111100000;
348:note_<=18'b100011000000000000;
349:note_<=18'b000011001111000000;
350:note_<=18'b100110000000000000;
351:note_<=18'b000110010110100000;
352:note_<=18'b100110000000000000;
353:note_<=18'b000110000111100000;
354:note_<=18'b100101000000000000;
355:note_<=18'b000101000111100000;
356:note_<=18'b100011000000000000;
357:note_<=18'b000011000111100000;
358:note_<=18'b100101000000000000;
359:note_<=18'b000101001111000000;
360:note_<=18'b100110000000000000;
361:note_<=18'b000110001111000000;
362:note_<=18'b101000000000000000;
363:note_<=18'b001000000111100000;
364:note_<=18'b100001000000000000;
365:note_<=18'b000001000111100000;
366:note_<=18'b100011000000000000;
367:note_<=18'b000011000111100000;
368:note_<=18'b100101000000000000;
369:note_<=18'b000101000111100000;
370:note_<=18'b100110000000000000;
371:note_<=18'b000110001111000000;
372:note_<=18'b101010000000000000;
373:note_<=18'b001010010110100000;
374:note_<=18'b101010000000000000;
375:note_<=18'b001010000111100000;
376:note_<=18'b101100000000000000;
377:note_<=18'b001100000111100000;
378:note_<=18'b101101000000000000;
379:note_<=18'b001101000111100000;
380:note_<=18'b110001000000000000;
381:note_<=18'b010001001111000000;
382:note_<=18'b101111000000000000;
383:note_<=18'b001111001111000000;
384:note_<=18'b101110000000000000;
385:note_<=18'b001110001111000000;
386:note_<=18'b101001000000000000;
387:note_<=18'b001001000111100000;
388:note_<=18'b101010000000000000;
389:note_<=18'b001010000111100000;
390:note_<=18'b101111000000000000;
391:note_<=18'b001111001111000000;
392:note_<=18'b101010000000000000;
393:note_<=18'b001010001111000000;
394:note_<=18'b101000000000000000;
395:note_<=18'b001000000111100000;
396:note_<=18'b110001000000000000;
397:note_<=18'b010001000111100000;
398:note_<=18'b101111000000000000;
399:note_<=18'b001111000111100000;
400:note_<=18'b101100000000000000;
401:note_<=18'b001100000111100000;
402:note_<=18'b101101000000000000;
403:note_<=18'b001101110100100000;
404:note_<=18'b101000000000000000;
405:note_<=18'b001000000011110000;
406:note_<=18'b100111000000000000;
407:note_<=18'b000111000011110000;
408:note_<=18'b101000000000000000;
409:note_<=18'b001000000111100000;
410:note_<=18'b100101000000000000;
411:note_<=18'b000101000111100000;
412:note_<=18'b100101000000000000;
413:note_<=18'b000101001011010000;
414:note_<=18'b100011000000000000;
415:note_<=18'b000011000011110000;
416:note_<=18'b100001000000000000;
417:note_<=18'b000001000111100000;
418:note_<=18'b100101000000000000;
419:note_<=18'b000101000111100000;
420:note_<=18'b100101000000000000;
421:note_<=18'b000101001111000000;
422:note_<=18'b100110000000000000;
423:note_<=18'b000110000011110000;
424:note_<=18'b100110000000000000;
425:note_<=18'b000110000011110000;
426:note_<=18'b100101000011110000;
427:note_<=18'b000101000011110000;
428:note_<=18'b100110000000000000;
429:note_<=18'b000110000001010001;
430:note_<=18'b101000000000000000;
431:note_<=18'b001000000000110011;
432:note_<=18'b101010000000000000;
433:note_<=18'b001010000000101000;
434:note_<=18'b100110000000000000;
435:note_<=18'b000110000001101001;
436:note_<=18'b100101000000000000;
437:note_<=18'b000101000000001001;
438:note_<=18'b100110000000000000;
439:note_<=18'b000110000010011001;
440:note_<=18'b100011000000000000;
441:note_<=18'b000011000000001111;
442:note_<=18'b100011000000000000;
443:note_<=18'b000011000000101111;
444:note_<=18'b100001000000000000;
445:note_<=18'b000001000010011001;
446:note_<=18'b100000000000000000;
447:note_<=18'b000000000001111010;
448:note_<=18'b100011000000000000;
449:note_<=18'b000011000001000000;
450:note_<=18'b100011000000000000;
451:note_<=18'b000011001110111101;
452:note_<=18'b100101000000000000;
453:note_<=18'b000101000011110000;
454:note_<=18'b100101000000000000;
455:note_<=18'b000101000011110000;
default: note_ <= 18'b0;
endcase

note_on <= note_[17:17];
note <= note_[16:12];
delay <= note_[11:0];
end
endmodule


