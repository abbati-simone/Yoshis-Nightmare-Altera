parameter ROMS_number=1;
parameter note_max_bits=5;
parameter address_max_bits=9;
parameter delay_max_bits=12;
parameter ticks_per_beat=960;
parameter BPM=84;
parameter BPS=1.4;
parameter ticks_hz=1344;
parameter delay_clocks_per_tick=1000;
parameter delay_clock_hz=1344000;
parameter delay_reg_bits=33;

