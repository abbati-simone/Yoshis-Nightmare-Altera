module notes_sequence_Yoshi_0(
	input clk,
	input [7:0] address,
	output reg [4:0] note,
	output reg note_on,
	output reg [9:0] delay
);

reg [15:0] note_;

always @(posedge clk) begin
case(address)
0:note_<=16'b1010011111000000;
1:note_<=16'b0010011001011000;
2:note_<=16'b1010000000000000;
3:note_<=16'b0010000001111000;
4:note_<=16'b1010010000000000;
5:note_<=16'b0010010001111000;
6:note_<=16'b1010100000000000;
7:note_<=16'b0010100001111000;
8:note_<=16'b1011000000000000;
9:note_<=16'b0011000101101000;
10:note_<=16'b1010010000000000;
11:note_<=16'b0010010001111000;
12:note_<=16'b1001010000000000;
13:note_<=16'b0001010001111000;
14:note_<=16'b1001000000000000;
15:note_<=16'b0001000001111000;
16:note_<=16'b1001010000000000;
17:note_<=16'b0001010001111000;
18:note_<=16'b1010010000000000;
19:note_<=16'b0010010001111000;
20:note_<=16'b1001110000000000;
21:note_<=16'b0001110011110000;
22:note_<=16'b1000100000000000;
23:note_<=16'b0000100011110000;
24:note_<=16'b1001110000000000;
25:note_<=16'b0001110011110000;
26:note_<=16'b1010010000000000;
27:note_<=16'b0010010011110000;
28:note_<=16'b1001110000000000;
29:note_<=16'b0001110111100000;
30:note_<=16'b1001010001111000;
31:note_<=16'b0001010001111000;
32:note_<=16'b1001000000000000;
33:note_<=16'b0001000001111000;
34:note_<=16'b1000100000000000;
35:note_<=16'b0000100001111000;
36:note_<=16'b1000000000000000;
37:note_<=16'b0000000101101000;
38:note_<=16'b1001110000000000;
39:note_<=16'b0001110001111000;
40:note_<=16'b1011000000000000;
41:note_<=16'b0011000011110000;
42:note_<=16'b1001110000000000;
43:note_<=16'b0001110011110000;
44:note_<=16'b1000000000000000;
45:note_<=16'b0000000101101000;
46:note_<=16'b1001110000000000;
47:note_<=16'b0001110001111000;
48:note_<=16'b1011000000000000;
49:note_<=16'b0011000011110000;
50:note_<=16'b1001110000000000;
51:note_<=16'b0001110011110000;
52:note_<=16'b1010010000000000;
53:note_<=16'b0010010011110000;
54:note_<=16'b1010010000000000;
55:note_<=16'b0010010010110100;
56:note_<=16'b1010010000000000;
57:note_<=16'b0010010000111100;
58:note_<=16'b1001110000000000;
59:note_<=16'b0001110001111000;
60:note_<=16'b1010010000000000;
61:note_<=16'b0010010001111000;
62:note_<=16'b1010100000000000;
63:note_<=16'b0010100001111000;
64:note_<=16'b1001110000000000;
65:note_<=16'b0001110001111000;
66:note_<=16'b1001010000000000;
67:note_<=16'b0001011001011000;
68:note_<=16'b1001010000000000;
69:note_<=16'b0001010001111000;
70:note_<=16'b1001110000000000;
71:note_<=16'b0001110001111000;
72:note_<=16'b1010010000000000;
73:note_<=16'b0010010001111000;
74:note_<=16'b1010100000000000;
75:note_<=16'b0010100011110000;
76:note_<=16'b1010100000000000;
77:note_<=16'b0010100011110000;
78:note_<=16'b1011100000000000;
79:note_<=16'b0011100011110000;
80:note_<=16'b1010100000000000;
81:note_<=16'b0010100011110000;
82:note_<=16'b1011000000000000;
83:note_<=16'b0011000001111000;
84:note_<=16'b1011000000000000;
85:note_<=16'b0011000011110000;
86:note_<=16'b1010100000000000;
87:note_<=16'b0010100001111000;
88:note_<=16'b1010010000000000;
89:note_<=16'b0010010111100000;
90:note_<=16'b1001110000000000;
91:note_<=16'b0001110001111000;
92:note_<=16'b1001110000000000;
93:note_<=16'b0001110011110000;
94:note_<=16'b1010010000000000;
95:note_<=16'b0010010001111000;
96:note_<=16'b1010110000000000;
97:note_<=16'b0010110011110000;
98:note_<=16'b1001110000000000;
99:note_<=16'b0001110011110000;
100:note_<=16'b1011000000000000;
101:note_<=16'b0011000001111000;
102:note_<=16'b1011000000000000;
103:note_<=16'b0011000011110000;
104:note_<=16'b1011100000000000;
105:note_<=16'b0011100001111000;
106:note_<=16'b1011000000000000;
107:note_<=16'b0011000001111000;
108:note_<=16'b1011000000000000;
109:note_<=16'b0011000001111000;
110:note_<=16'b1011100000000000;
111:note_<=16'b0011100001111000;
112:note_<=16'b1100000000000000;
113:note_<=16'b0100000001111000;
114:note_<=16'b1100010000000000;
115:note_<=16'b0100010111100000;
116:note_<=16'b1011000000000000;
117:note_<=16'b0011000111100000;
118:note_<=16'b1011100000000000;
119:note_<=16'b0011100001111000;
120:note_<=16'b1011100000000000;
121:note_<=16'b0011100011110000;
122:note_<=16'b1100000000000000;
123:note_<=16'b0100000001111000;
124:note_<=16'b1100010000000000;
125:note_<=16'b0100010011110000;
126:note_<=16'b1011100000000000;
127:note_<=16'b0011100011110000;
128:note_<=16'b1011000000000000;
129:note_<=16'b0011000010110100;
130:note_<=16'b1011100000000000;
131:note_<=16'b0011100000111100;
132:note_<=16'b1011000000000000;
133:note_<=16'b0011000001111000;
134:note_<=16'b1011100000000000;
135:note_<=16'b0011100001111000;
136:note_<=16'b1011000000000000;
137:note_<=16'b0011000001111000;
138:note_<=16'b1010100000000000;
139:note_<=16'b0010100001111000;
140:note_<=16'b1010010000000000;
141:note_<=16'b0010010001111000;
142:note_<=16'b1001110000000000;
143:note_<=16'b0001110001111000;
144:note_<=16'b1001010000000000;
145:note_<=16'b0001010111100000;
default: note_ <= 16'b0;
endcase

note_on <= note_[15:15];
note <= note_[14:10];
delay <= note_[9:0];
end
endmodule


