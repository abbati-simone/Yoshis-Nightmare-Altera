parameter ROM_0_messages_len=456;
parameter ROM_0_note_min=66;
parameter ROM_0_note_max=83;
parameter ROM_0_delay_min=0;
parameter ROM_0_delay_max=3360;
parameter ROM_0_messages_address_bits=9;
parameter ROM_0_note_nbit=5;
parameter ROM_0_delay_nbit=12;

